library verilog;
use verilog.vl_types.all;
entity SLC3_2 is
end SLC3_2;
