library verilog;
use verilog.vl_types.all;
entity test_memory_sv_unit is
end test_memory_sv_unit;
